netcdf hycom1_75 {
dimensions:
	layers = 75 ;
	interfaces = 76 ;
variables:
	double dz(layers) ;
		dz:long_name = "z* coordinate level thickness" ;
		dz:units = "m" ;
	double sigma2(interfaces) ;
		sigma2:long_name = "Interface target potential density referenced to 2000 dbars" ;
		sigma2:units = "kg/m3" ;
data:

 dz = 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2.01, 2.01, 2.02, 2.03, 2.04, 2.06, 
    2.08, 2.12, 2.16, 2.22, 2.3, 2.4, 2.52, 2.67, 2.85, 3.08, 3.35, 3.68, 
    4.08, 4.54, 5.1, 5.75, 6.51, 7.39, 8.42, 9.6, 10.96, 12.51, 14.28, 16.3, 
    18.58, 21.16, 24.07, 27.33, 30.99, 35.07, 39.63, 44.69, 50.32, 56.54, 
    63.42, 71.01, 79.37, 88.55, 98.63, 109.66, 121.72, 134.89, 149.24, 
    164.86, 181.84, 200.27, 220.25, 241.88, 265.27, 290.52, 317.76, 347.12, 
    378.71, 412.68, 449.16, 488.31, 530.27, 575.19 ;

 sigma2 = 1010, 1014.3034, 1017.8088, 1020.843, 1023.5566, 1025.813, 
    1027.0275, 1027.9114, 1028.6422, 1029.2795, 1029.852, 1030.3762, 
    1030.8626, 1031.3183, 1031.7486, 1032.1572, 1032.5471, 1032.9207, 
    1033.2798, 1033.6261, 1033.9608, 1034.2519, 1034.4817, 1034.6774, 
    1034.8508, 1035.0082, 1035.1533, 1035.2886, 1035.4159, 1035.5364, 
    1035.6511, 1035.7608, 1035.8661, 1035.9675, 1036.0645, 1036.1554, 
    1036.2411, 1036.3223, 1036.3998, 1036.4739, 1036.5451, 1036.6137, 
    1036.68, 1036.7441, 1036.8062, 1036.8526, 1036.8874, 1036.9164, 
    1036.9418, 1036.9647, 1036.9857, 1037.0052, 1037.0236, 1037.0409, 
    1037.0574, 1037.0738, 1037.0902, 1037.1066, 1037.123, 1037.1394, 
    1037.1558, 1037.1722, 1037.1887, 1037.206, 1037.2241, 1037.2435, 
    1037.2642, 1037.2866, 1037.3112, 1037.3389, 1037.3713, 1037.4118, 
    1037.475, 1037.6332, 1037.8104, 1038 ;
}
