../../OM4_025/INPUT/hycom1_75.cdl