../../common_BML/zgrid.cdl