../../OM4_025/INPUT/hycom1_75_800m.cdl