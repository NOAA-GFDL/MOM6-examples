netcdf hycom1_50 {
dimensions:
	layers = 50 ;
	interfaces = 51 ;
variables:
	double dz(layers) ;
		dz:long_name = "z* coordinate level thickness" ;
		dz:units = "m" ;
	double sigma2(interfaces) ;
		sigma2:long_name = "Interface target potential density referenced to 2000 dbars" ;
		sigma2:units = "kg/m3" ;
data:

 dz = 5, 5, 5, 5, 5.1, 5.2, 5.3, 5.4, 5.5, 6, 7, 8, 
    9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 
    21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30 ;

 sigma2 = 1010, 1016.1289, 1020.843, 1024.821, 1027.0275, 1028.2911, 
    1029.2795, 1030.1194, 1030.8626, 1031.5364, 1032.1572, 1032.7358, 
    1033.2798, 1033.7948, 1034.2519, 1034.5828, 1034.8508, 1035.0821, 
    1035.2886, 1035.4769, 1035.6511, 1035.814, 1035.9675, 1036.1107, 
    1036.2411, 1036.3615, 1036.4739, 1036.5797, 1036.68, 1036.7755, 
    1036.8526, 1036.9024, 1036.9418, 1036.9754, 1037.0052, 1037.0323, 
    1037.0574, 1037.082, 1037.1066, 1037.1312, 1037.1558, 1037.1804, 
    1037.206, 1037.2337, 1037.2642, 1037.2986, 1037.3389, 1037.3901, 
    1037.475, 1037.7204, 1038 ;
}
