netcdf interface_IC_2layer {
dimensions:
        nki = 3 ; // (47 currently)
variables:
        double eta(nki) ;
                eta:long_name = "Initial depth of interfaces" ;
                eta:units = "meters" ;
data:

 eta = 0, -700., -12000. ;

}
