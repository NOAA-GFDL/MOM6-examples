netcdf zgrid {
dimensions:
	zt = 35 ;
	zw = 36 ;
variables:
	double zt(zt) ;
		zt:long_name = "Diagnostic depth coordinate layer position" ;
		zt:comment = "Used for diagnostics only." ;
		zt:units = "m" ;
	double zw(zw) ;
		zw:long_name = "Diagnostic depth coordinate interface position" ;
		zw:comment = "Used for diagnostics only." ;
		zw:units = "m" ;

// global attributes:
		:filename = "vgrid_75_2m.nc" ;
data:

 zt = 0.5, 1.5, 2.5, 3.5, 5, 7, 9, 11, 13, 15, 17, 19, 22.5, 27.5, 32.5, 
    37.5, 42.5, 47.5, 55, 65, 75, 85, 95, 110, 130, 150, 170, 190, 210, 230, 
    250, 270, 290, 325, 375 ;

 zw = 0, 1, 2, 3, 4, 6, 8, 10, 12, 14, 16, 18, 20, 25, 30, 35, 40, 45, 50, 
    60, 70, 80, 90, 100, 120, 140, 160, 180, 200, 220, 240, 260, 280, 300, 
    350, 400 ;
}
