netcdf vgrid_75_2m_575m {
dimensions:
	nz = 75 ;
variables:
	double dz(nz) ;
		dz:long_name = "z* coordinate level thickness" ;
		dz:units = "m" ;

// global attributes:
		:filename = "vgrid_75_2m_575m.nc" ;
data:

 dz = 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2.01, 2.01, 2.02, 2.03, 2.04, 2.06, 
    2.08, 2.12, 2.16, 2.22, 2.3, 2.4, 2.52, 2.67, 2.85, 3.08, 3.35, 3.68, 
    4.08, 4.54, 5.1, 5.75, 6.51, 7.39, 8.42, 9.6, 10.96, 12.51, 14.28, 16.3, 
    18.58, 21.16, 24.07, 27.33, 30.99, 35.07, 39.63, 44.69, 50.32, 56.54, 
    63.42, 71.01, 79.37, 88.55, 98.63, 109.66, 121.72, 134.89, 149.24, 
    164.86, 181.84, 200.27, 220.25, 241.88, 265.27, 290.52, 317.76, 347.12, 
    378.71, 412.68, 449.16, 488.31, 530.27, 575.19 ;
}
