../../OM4_05/INPUT/analysis_vgrid_lev35.v1.cdl