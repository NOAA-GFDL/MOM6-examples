netcdf zgrid {
dimensions:
	zt = 60 ;
	zw = 61 ;
variables:
	double zt(zt) ;
		zt:long_name = "Depth of Level Center" ;
		zt:units = "m" ;
		zt:positive = "down" ;
	double zw(zw) ;
		zw:long_name = "Depth of edges" ;
		zw:units = "m" ;
		zw:positive = "down" ;

// global attributes:
		:filename = "zgrid.nc" ;
data:

 zt = 5, 15, 25, 35, 45, 55, 65, 75, 85, 95, 105, 115, 125, 135, 145, 155, 
    165, 175, 185, 195, 205, 215, 225, 235, 245, 255, 265, 275, 285, 295, 
    305, 315, 325, 335, 345, 355, 365, 375, 385, 395, 405, 415, 425, 435, 
    445, 455, 465, 475, 485, 495, 510, 530, 550, 570, 590, 625, 675, 725, 
    775, 850 ;

 zw = 0, 10, 20, 30, 40, 50, 60, 70, 80, 90, 100, 110, 120, 130, 140, 150, 
    160, 170, 180, 190, 200, 210, 220, 230, 240, 250, 260, 270, 280, 290, 
    300, 310, 320, 330, 340, 350, 360, 370, 380, 390, 400, 410, 420, 430, 
    440, 450, 460, 470, 480, 490, 500, 520, 540, 560, 580, 600, 650, 700, 
    750, 800, 900 ;
}
