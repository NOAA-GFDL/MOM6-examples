../../common_EPBL/zgrid.cdl