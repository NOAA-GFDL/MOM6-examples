netcdf diag_rho2 {
dimensions:
	Interface = 65 ;
variables:
	double rho2(Interface) ;
		rho2:units = "kg m-3" ;
data:

 rho2 = 997, 1011.4925, 1015.6375, 1019.7825, 1023.9275, 1028.0725, 1030.591, 
    1031.378, 1031.974, 1032.431, 1032.8055, 1033.133, 1033.4315, 1033.7105, 
    1033.9745, 1034.225, 1034.462, 1034.685, 1034.894, 1035.088, 1035.2665, 
    1035.4295, 1035.5775, 1035.712, 1035.8335, 1035.9435, 1036.044, 
    1036.1365, 1036.222, 1036.302, 1036.378, 1036.451, 1036.522, 1036.591, 
    1036.659, 1036.725, 1036.7855, 1036.8385, 1036.884, 1036.924, 1036.959, 
    1036.989, 1037.015, 1037.0375, 1037.0575, 1037.0755, 1037.092, 1037.108, 
    1037.124, 1037.14, 1037.156, 1037.172, 1037.188, 1037.205, 1037.224, 
    1037.246, 1037.274, 1037.315, 1037.375, 1037.455, 1037.56, 1037.69, 
    1037.83, 1037.97, 1039 ;
}
