netcdf vgrid_75_2m {
dimensions:
	nz = 75 ;
variables:
	double dz(nz) ;
		dz:long_name = "z coordinate level thickness" ;
		dz:units = "m" ;

// global attributes:
		:filename = "vgrid_75_2m.nc" ;
data:

 dz = 2, 2, 2, 2, 2.01, 2.01, 2.02, 2.03, 2.05, 2.08, 2.11, 2.15, 2.2, 2.27, 
    2.34, 2.44, 2.55, 2.69, 2.85, 3.04, 3.27, 3.54, 3.85, 4.22, 4.66, 5.18, 
    5.79, 6.52, 7.37, 8.37, 9.55, 10.94, 12.57, 14.48, 16.72, 19.33, 22.36, 
    25.87, 29.91, 34.53, 39.79, 45.72, 52.37, 59.76, 67.89, 76.74, 86.29, 
    96.47, 107.2, 118.35, 129.81, 141.42, 153.01, 164.41, 175.47, 186.01, 
    195.9, 205.01, 213.27, 220.6, 226.99, 232.43, 236.96, 240.63, 243.52, 
    245.72, 247.33, 248.45, 249.18, 249.62, 249.86, 249.96, 249.99, 250, 250 ;
}
