../../OM4_05/INPUT/hycom1_75_800m.cdl