../../OM4_025/INPUT/vgrid_75_2m.cdl