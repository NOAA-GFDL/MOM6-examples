netcdf vgrid {
dimensions:
	nk = 80 ;
	nkp1 = 81 ;
variables:
	double dz(nk) ;
		dz:long_name = "z coordinate level thickness" ;
		dz:units = "m" ;
	double zt(nk) ;
		zt:long_name = "Diagnostic z coordinate level position" ;
		zt:comment = "Used for diagnostics only" ;
		zt:units = "m" ;
	double zw(nkp1) ;
		zw:long_name = "Diagnostic z coordinate interface position" ;
		zw:comment = "Used for diagnostics only" ;
		zw:units = "m" ;

// global attributes:
		:filename = "vgrid.nc" ;
data:

 dz = 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 
      2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 
      2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 
      2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 
      5., 5., 5., 5., 5., 5., 5., 5., 5., 5., 
      5., 5., 5., 5., 5., 5., 5., 5., 5., 5.,
      10., 10., 10., 10., 10., 10., 10., 10., 10., 10.,  
      100.,100.,250.,250.,500.,500.,500.,500.,500.,500. ;

 zt = 1.25,3.75,6.25,8.75,11.25,13.75,16.25,18.75,21.25,23.75,
      26.25,28.75,31.25,33.75,36.25,38.75,41.25,43.75,46.25,48.75,
      51.25,53.75,56.25,58.75,61.25,63.75,66.25,68.75,71.25,73.75,
      76.25,78.75,81.25,83.75,86.25,88.75,91.25,93.75,96.25,98.75,
      102.5,107.5,112.5,117.5,122.5,127.5,132.5,137.5,142.5,147.5,
      152.5,157.5,162.5,167.5,172.5,177.5,182.5,187.5,192.5,197.5,
      205.,215.,225.,235.,245.,255.,265.,275.,285.,295.,
      350.,450.,625.,875.,1250.,1750.,2250.,2750.,3250.,3750. ;

 zw = 0.,2.5,5.,7.5,10.,12.5,15.,17.5,20.,22.5,25.,
      27.5,30.,32.5,35.,37.5,40.,42.5,45.,47.5,50.,
      50.,52.5,55.,57.5,60.,62.5,65.,67.5,70.,72.5,75.,
      77.5,80.,82.5,85.,87.5,90.,92.5,95.,97.5,100.,
      105.,110.,115.,120.,125.,130.,135.,140.,145.,150.,
      155.,160.,165.,170.,175.,180.,185.,190.,195.,200.,
      210.,220.,230.,240.,250.,260.,270.,280.,290.,300.,
      400.,500.,750.,1000.,1500.,2000.,2500.,3000.,3500.,4000. ;
      
}
