../../common_KPP/zgrid.cdl